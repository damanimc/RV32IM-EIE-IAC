module DataMem#(
  parameter DATA_WIDTH = 32

)(
input logic clk,
input logic [DATA_WIDTH-1:0] a,
input logic [2:0] memCtrl,
input logic we,
input logic [DATA_WIDTH-1:0] wd,
output logic[DATA_WIDTH-1:0] rd
);

logic [7:0] ram_array [20'h1FFFF:0];//byte addressable up to where the data memory goes

// initial begin
//     $readmemh("sinerom.mem", rom_array);
// end;

//can take out wd3 enable in alutop/ 
//always_comb for asynchronous logi
assign rd = {ram_array[a+3], ram_array[a+2], ram_array[a+1], ram_array[a]};//whole word

//passing unaligned address 
initial begin 
    $display("Loading RAM...");
    $readmemh("Data.mem",ram_array,20'h10000);
end;

always_comb //load
case(memCtrl[2])
  1'b0:begin

    case(memCtrl[1:0])
      2'b00: rd= {{24{ram_array[a][7]}},ram_array[a]};
      2'b01: rd= {{16{ram_array[a+1][7]}},ram_array[a+1], ram_array[a]};
      2'b10: rd= {ram_array[a+3], ram_array[a+2], ram_array[a+1], ram_array[a]};
    endcase 
  end
  1'b1:begin //zero extend
    case(memCtrl[1:0])
    2'b00: rd= {24'b0,ram_array[a]};
    2'b01: rd= {16'b0,ram_array[a+1], ram_array[a]};
    endcase
  end 
endcase


 
always_ff @(posedge clk) //store 
if(we)
  case(memCtrl[1:0])
            2'b00: ram_array[a] <= wd[7:0];
            2'b01: {ram_array[a+1], ram_array[a]}<=wd[15:0];
            2'b10: {ram_array[a+3], ram_array[a+2], ram_array[a+1], ram_array[a]}<=wd[31:0];
  endcase 
endmodule

